library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.MyPackage.all;
entity DEC32 is
    Port ( sel : in  STD_LOGIC_VECTOR (4 downto 0);
           o : out  STD_LOGIC_VECTOR (31 downto 0));
end DEC32;

architecture Behavioral of DEC32 is

begin

o<="00000000000000000000000000000001" when sel= "00000" else
	"00000000000000000000000000000010" when sel= "00001" else
	"00000000000000000000000000000100" when sel= "00010" else
	"00000000000000000000000000001000" when sel= "00011" else
	"00000000000000000000000000010000" when sel= "00100" else
	"00000000000000000000000000100000" when sel= "00101" else
	"00000000000000000000000001000000" when sel= "00110" else
	"00000000000000000000000010000000" when sel= "00111" else
	"00000000000000000000000100000000" when sel= "01000" else
	"00000000000000000000001000000000" when sel= "01001" else
	"00000000000000000000010000000000" when sel= "01010" else
	"00000000000000000000100000000000" when sel= "01011" else
	"00000000000000000001000000000000" when sel= "01100" else
	"00000000000000000010000000000000" when sel= "01101" else
	"00000000000000000100000000000000" when sel= "01110" else
	"00000000000000001000000000000000" when sel= "01111" else
	"00000000000000010000000000000000" when sel= "10000" else
	"00000000000000100000000000000000" when sel= "10001" else
	"00000000000001000000000000000000" when sel= "10010" else
	"00000000000010000000000000000000" when sel= "10011" else
	"00000000000100000000000000000000" when sel= "10100" else
	"00000000001000000000000000000000" when sel= "10101" else
	"00000000010000000000000000000000" when sel= "10110" else
	"00000000100000000000000000000000" when sel= "10111" else
	"00000001000000000000000000000000" when sel= "11000" else
	"00000010000000000000000000000000" when sel= "11001" else
	"00000100000000000000000000000000" when sel= "11010" else
	"00001000000000000000000000000000" when sel= "11011" else
	"00010000000000000000000000000000" when sel= "11100" else
	"00100000000000000000000000000000" when sel= "11101" else
	"01000000000000000000000000000000" when sel= "11110" else
	"10000000000000000000000000000000" when sel= "11111" ;
end Behavioral;

